* C:\Users\Petter\Documents\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Fri Sep 21 15:41:01 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
