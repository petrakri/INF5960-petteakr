* C:\Users\Petter\Documents\prog\github\INF5960-petteakr\pspice\Schematics\inverting_opamp.sch

* Schematics Version 9.1 - Web Update 1
* Tue Mar 05 16:02:20 2019



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "inverting_opamp.net"
.INC "inverting_opamp.als"


.probe


.END
