* C:\Users\Petter\Documents\prog\github\INF5960-petteakr\pspice\Schematics\noninvertin_opamp.sch

* Schematics Version 9.1 - Web Update 1
* Fri Oct 12 15:06:51 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "noninvertin_opamp.net"
.INC "noninvertin_opamp.als"


.probe


.END
